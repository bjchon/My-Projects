** Profile: "SCHEMATIC1-sim2"  [ c:\users\bdawg\onedrive\desktop\uc merced\summer 2022\engr 065 circuit theory\lab\lab9\2\lab9circuit2-PSpiceFiles\SCHEMATIC1\sim2.sim ] 

** Creating circuit file "sim2.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 2ms 0 5us 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
